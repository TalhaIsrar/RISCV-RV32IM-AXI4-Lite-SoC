module led(
    input clk,
    input rst,
    input [7:0] led_write
);
    

endmodule